module tb_freq_div;




endmodule
