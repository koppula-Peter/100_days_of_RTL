module tb_shift_reg;




endmodule
