module tb_overflow;
  
