module tb_clock_generator;

  
