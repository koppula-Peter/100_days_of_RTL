moduel shift_reg(input in, output reg out);




endmodule
