module freq_divider(input freq_in,index,rst,output freq_out);


endmodule
